module jaltop #(
    parameter WIDTH = 32

)(

   input logic [2:0] PCSrc,
   input logic ALUResult
);

    

