`ifndef DEF_SV

    `define DEF_SV
    `define PC_NEXT                 3'b000
    `define PC_ALWAYS               3'b001
    `define PC_JALR                 3'b010
    `define PC_INV_COND             3'b100
    `define PC_COND                 3'b101

`endif