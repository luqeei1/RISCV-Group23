`ifndef DEF_SV

    `define DEF_SV

    `define PC_NEXT                 2'b00
    `define PC_JUMP                 2'b01
    `define PC_JALR                 2'b11
    `define PC_COND_JUMP            2'b10

`endif
