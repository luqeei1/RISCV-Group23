// add once done
