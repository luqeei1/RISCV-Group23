module instructionMemory #(
    parameter ADDRESS_WIDTH = 32,
              DATA_WIDTH = 32
)(
    input logic [31:0]                  PC,
    output logic [DATA_WIDTH-1:0] instr
);

logic [7:0] rom_array [2**16 - 1 : 0];


initial begin
    $display("Loading rom.");
    $readmemh("program.hex", rom_array);     
    $display("ROM loaded successfully.");
end

// Check if PC is in the valid range

// Fetch instruction only if address is valid, 0 otherwise
assign instr = {{rom_array[PC + 3]}, {rom_array[PC + 2]}, {rom_array[PC + 1]}, {rom_array[PC]}};

endmodule
